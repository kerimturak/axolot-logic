module tb_ders_001();
    wire a;
    wire b;

    ders_001 uut (
        .a(a),
        .b(b)
    );
endmodule