module ders_002(
    input a,
    output b
);
    assign b = a;
endmodule