module ders_001 (
    input  a,
    output b
);
  assign b = a;
endmodule
